PACKAGE common IS
    TYPE state IS (START, STOP, READ, WRITE, IDLE, DONE, SEND, RCV);
END common;