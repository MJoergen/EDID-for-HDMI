LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE dataBytes IS
    TYPE data IS ARRAY (1 TO 256) OF STD_LOGIC_VECTOR (7 DOWNTO 0);
END PACKAGE;
